///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: SameBit
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbench();
`include "../Test/Test.v"
///////////////////////////////////////////////////////////////////////////////////
// Input: A (1-bit)
reg A;
///////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////
// Output: S (1-bit)
wire S;
///////////////////////////////////////////////////////////////////////////////////

SameBit mySame(.Ain(A), .Aout(S));

initial begin
////////////////////////////////////////////////////////////////////////////////////////
// Test: A=0
$display("Testing: A=0");
A=0;   #10; 
verifyEqual(S, A);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: A=1
$display("Testing: A=1");
A=1;   #10; 
verifyEqual(S, A);
////////////////////////////////////////////////////////////////////////////////////////
$display("All tests passed.");
end

endmodule
